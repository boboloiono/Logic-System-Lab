`timescale 1ns/1ps
module problem2 (input d, input clk, output q, output q_bar);
endmodule