module problem3 (input d, input clk, output q, output q_bar);
endmodule