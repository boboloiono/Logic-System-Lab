module problem1 (input d, input c, output q, output q_bar);
endmodule